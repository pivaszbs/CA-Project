library verilog;
use verilog.vl_types.all;
entity simple_ram_tb is
    port(
        abidna          : out    vl_logic
    );
end simple_ram_tb;
