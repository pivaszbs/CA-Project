module rate_tb(output a);
	
	reg [31:0] data;
	reg [31:0] addr;
	reg wr;
	reg clk;
	reg state;
	wire is_missrate;
	reg[31:0] missrate_counter;
	reg[31:0] hitrate_counter;
	
	wire [31:0] out;
	
	cache_4way cache_4way(
	.data(data),
	.addr(addr),
	.wr(wr),	
	.clk(clk),
	.is_missrate(is_missrate),
	.out(out));
	
	reg init_state;
		
	initial
	begin
		init_state = 1;
		clk = 1;		
		state = 0;
		missrate_counter = 0;
		hitrate_counter = 0;
			
		data = 32'b00000000000000000000000000000001;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000010;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000011;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000100;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000101;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000110;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000000111;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001000;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001001;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001010;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001011;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001100;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001101;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001110;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000001111;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010000;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010001;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010010;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010011;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010100;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010101;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000010110;
addr = 32'b00000000000000000000011001110010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000000010111;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011000;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011001;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011010;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011011;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011100;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011101;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011110;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000011111;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100000;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100001;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100010;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100011;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100100;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100101;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100110;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000100111;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101000;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101001;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101010;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101011;
addr = 32'b00000000000000000000011001000101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000000101100;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101101;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101110;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000101111;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110000;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110001;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110010;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110011;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110100;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110101;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110110;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000110111;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111000;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111001;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111010;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111011;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111100;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111101;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111110;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000000111111;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000000;
addr = 32'b00000000000000000000011000011000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000001000001;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000010;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000011;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000100;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000101;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000110;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001000111;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001000;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001001;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001010;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001011;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001100;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001101;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001110;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001001111;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010000;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010001;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010010;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010011;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010100;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010101;
addr = 32'b00000000000000000000010111101011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000001010110;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001010111;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011000;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011001;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011010;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011011;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011100;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011101;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011110;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001011111;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100000;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100001;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100010;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100011;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100100;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100101;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100110;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001100111;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101000;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101001;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101010;
addr = 32'b00000000000000000000010110111110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000001101011;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101100;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101101;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101110;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001101111;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110000;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110001;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110010;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110011;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110100;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110101;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110110;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001110111;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111000;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111001;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111010;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111011;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111100;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111101;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111110;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000001111111;
addr = 32'b00000000000000000000010110010001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000010000000;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000001;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000010;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000011;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000100;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000101;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000110;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010000111;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001000;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001001;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001010;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001011;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001100;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001101;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001110;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010001111;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010000;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010001;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010010;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010011;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010100;
addr = 32'b00000000000000000000010101100100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000010010101;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010110;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010010111;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011000;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011001;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011010;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011011;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011100;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011101;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011110;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010011111;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100000;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100001;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100010;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100011;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100100;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100101;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100110;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010100111;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101000;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101001;
addr = 32'b00000000000000000000010100110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000010101010;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101011;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101100;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101101;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101110;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010101111;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110000;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110001;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110010;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110011;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110100;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110101;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110110;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010110111;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111000;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111001;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111010;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111011;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111100;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111101;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000010111110;
addr = 32'b00000000000000000000010100001010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000010111111;
addr = 32'b00000000000000000000000000000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000000;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000001;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000010;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000011;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000100;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000101;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000110;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011000111;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001000;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001001;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001010;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001011;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001100;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001101;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001110;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011001111;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010000;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010001;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010010;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010011;
addr = 32'b00000000000000000000010011011101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000011010100;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010101;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010110;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011010111;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011000;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011001;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011010;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011011;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011100;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011101;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011110;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011011111;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100000;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100001;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100010;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100011;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100100;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100101;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100110;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011100111;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101000;
addr = 32'b00000000000000000001101111101110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000011101001;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101010;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101011;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101100;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101101;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101110;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011101111;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110000;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110001;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110010;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110011;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110100;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110101;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110110;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011110111;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111000;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111001;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111010;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111011;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111100;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111101;
addr = 32'b00000000000000000001101101011101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000011111110;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000011111111;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000000;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000001;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000010;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000011;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000100;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000101;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000110;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100000111;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001000;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001001;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001010;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001011;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001100;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001101;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001110;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100001111;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010000;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010001;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010010;
addr = 32'b00000000000000000001101011001100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000100010011;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010100;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010101;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010110;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100010111;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011000;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011001;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011010;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011011;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011100;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011101;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011110;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100011111;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100000;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100001;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100010;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100011;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100100;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100101;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100110;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100100111;
addr = 32'b00000000000000000001101000111011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000100101000;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101001;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101010;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101011;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101100;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101101;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101110;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100101111;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110000;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110001;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110010;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110011;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110100;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110101;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110110;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100110111;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111000;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111001;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111010;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111011;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111100;
addr = 32'b00000000000000000001100110101010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000100111101;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111110;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000100111111;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000000;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000001;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000010;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000011;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000100;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000101;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000110;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101000111;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001000;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001001;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001010;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001011;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001100;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001101;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001110;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101001111;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010000;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010001;
addr = 32'b00000000000000000001100100011001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000101010010;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010011;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010100;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010101;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010110;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101010111;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011000;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011001;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011010;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011011;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011100;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011101;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011110;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101011111;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100000;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100001;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100010;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100011;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100100;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100101;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101100110;
addr = 32'b00000000000000000001100010001000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000101100111;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101000;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101001;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101010;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101011;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101100;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101101;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101110;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101101111;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110000;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110001;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110010;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110011;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110100;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110101;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110110;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101110111;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111000;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111001;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111010;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111011;
addr = 32'b00000000000000000001011111110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000101111100;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111101;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111110;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000101111111;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000000;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000001;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000010;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000011;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000100;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000101;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000110;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110000111;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001000;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001001;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001010;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001011;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001100;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001101;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001110;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110001111;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010000;
addr = 32'b00000000000000000001011101100110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000110010001;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010010;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010011;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010100;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010101;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010110;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110010111;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011000;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011001;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011010;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011011;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011100;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011101;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011110;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110011111;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100000;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100001;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100010;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100011;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100100;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100101;
addr = 32'b00000000000000000001011011010101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000110100110;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110100111;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101000;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101001;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101010;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101011;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101100;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101101;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101110;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110101111;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110000;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110001;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110010;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110011;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110100;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110101;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110110;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110110111;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111000;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111001;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111010;
addr = 32'b00000000000000000011000101101010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000110111011;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111100;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111101;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111110;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000110111111;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000000;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000001;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000010;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000011;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000100;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000101;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000110;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111000111;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001000;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001001;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001010;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001011;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001100;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001101;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001110;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111001111;
addr = 32'b00000000000000000011000001110101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000111010000;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010001;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010010;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010011;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010100;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010101;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010110;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111010111;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011000;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011001;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011010;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011011;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011100;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011101;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011110;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111011111;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100000;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100001;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100010;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100011;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100100;
addr = 32'b00000000000000000010111110000000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000111100101;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100110;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111100111;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101000;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101001;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101010;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101011;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101100;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101101;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101110;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111101111;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110000;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110001;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110010;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110011;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110100;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110101;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110110;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111110111;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111000;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111001;
addr = 32'b00000000000000000010111010001011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000000111111010;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111011;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111100;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111101;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111110;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000000111111111;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000000;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000001;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000010;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000011;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000100;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000101;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000110;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000000111;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001000;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001001;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001010;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001011;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001100;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001101;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000001110;
addr = 32'b00000000000000000010110110010110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001000001111;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010000;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010001;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010010;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010011;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010100;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010101;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010110;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000010111;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011000;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011001;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011010;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011011;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011100;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011101;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011110;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000011111;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100000;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100001;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100010;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100011;
addr = 32'b00000000000000000010110010100001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001000100100;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100101;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100110;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000100111;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101000;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101001;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101010;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101011;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101100;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101101;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101110;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000101111;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110000;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110001;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110010;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110011;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110100;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110101;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110110;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000110111;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111000;
addr = 32'b00000000000000000010101110101100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001000111001;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111010;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111011;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111100;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111101;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111110;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001000111111;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000000;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000001;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000010;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000011;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000100;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000101;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000110;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001000111;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001000;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001001;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001010;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001011;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001100;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001101;
addr = 32'b00000000000000000010101010110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001001001110;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001001111;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010000;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010001;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010010;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010011;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010100;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010101;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010110;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001010111;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011000;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011001;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011010;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011011;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011100;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011101;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011110;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001011111;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100000;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100001;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100010;
addr = 32'b00000000000000000010100111000010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001001100011;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100100;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100101;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100110;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001100111;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101000;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101001;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101010;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101011;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101100;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101101;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101110;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001101111;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110000;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110001;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110010;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110011;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110100;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110101;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110110;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001110111;
addr = 32'b00000000000000000010100011001101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001001111000;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111001;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111010;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111011;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111100;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111101;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111110;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001001111111;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000000;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000001;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000010;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000011;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000100;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000101;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000110;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010000111;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001000;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001001;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001010;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001011;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001100;
addr = 32'b00000000000000000100011011100110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001010001101;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001110;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010001111;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010000;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010001;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010010;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010011;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010100;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010101;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010110;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010010111;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011000;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011001;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011010;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011011;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011100;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011101;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011110;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010011111;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100000;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100001;
addr = 32'b00000000000000000100010110001101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001010100010;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100011;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100100;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100101;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100110;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010100111;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101000;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101001;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101010;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101011;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101100;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101101;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101110;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010101111;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110000;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110001;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110010;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110011;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110100;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110101;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010110110;
addr = 32'b00000000000000000100010000110100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001010110111;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111000;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111001;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111010;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111011;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111100;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111101;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111110;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001010111111;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000000;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000001;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000010;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000011;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000100;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000101;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000110;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011000111;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001000;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001001;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001010;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001011;
addr = 32'b00000000000000000100001011011011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001011001100;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001101;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001110;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011001111;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010000;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010001;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010010;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010011;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010100;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010101;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010110;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011010111;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011000;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011001;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011010;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011011;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011100;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011101;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011110;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011011111;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100000;
addr = 32'b00000000000000000100000110000010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001011100001;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100010;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100011;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100100;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100101;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100110;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011100111;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101000;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101001;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101010;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101011;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101100;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101101;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101110;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011101111;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110000;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110001;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110010;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110011;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110100;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110101;
addr = 32'b00000000000000000100000000101001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001011110110;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011110111;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111000;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111001;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111010;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111011;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111100;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111101;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111110;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001011111111;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000000;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000001;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000010;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000011;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000100;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000101;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000110;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100000111;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001000;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001001;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001010;
addr = 32'b00000000000000000011111011010000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001100001011;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001100;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001101;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001110;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100001111;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010000;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010001;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010010;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010011;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010100;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010101;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010110;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100010111;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011000;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011001;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011010;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011011;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011100;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011101;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011110;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100011111;
addr = 32'b00000000000000000011110101110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001100100000;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100001;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100010;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100011;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100100;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100101;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100110;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100100111;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101000;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101001;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101010;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101011;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101100;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101101;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101110;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100101111;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110000;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110001;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110010;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110011;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110100;
addr = 32'b00000000000000000011110000011110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001100110101;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110110;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100110111;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111000;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111001;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111010;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111011;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111100;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111101;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111110;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001100111111;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000000;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000001;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000010;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000011;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000100;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000101;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000110;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101000111;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001000;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001001;
addr = 32'b00000000000000000011101011000101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001101001010;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001011;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001100;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001101;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001110;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101001111;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010000;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010001;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010010;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010011;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010100;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010101;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010110;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101010111;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011000;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011001;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011010;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011011;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011100;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011101;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101011110;
addr = 32'b00000000000000000101110001100010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001101011111;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100000;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100001;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100010;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100011;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100100;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100101;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100110;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101100111;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101000;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101001;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101010;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101011;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101100;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101101;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101110;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101101111;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110000;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110001;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110010;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110011;
addr = 32'b00000000000000000101101010100101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001101110100;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110101;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110110;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101110111;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111000;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111001;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111010;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111011;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111100;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111101;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111110;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001101111111;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000000;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000001;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000010;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000011;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000100;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000101;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000110;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110000111;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001000;
addr = 32'b00000000000000000101100011101000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001110001001;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001010;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001011;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001100;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001101;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001110;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110001111;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010000;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010001;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010010;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010011;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010100;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010101;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010110;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110010111;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011000;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011001;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011010;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011011;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011100;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011101;
addr = 32'b00000000000000000101011100101011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001110011110;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110011111;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100000;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100001;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100010;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100011;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100100;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100101;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100110;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110100111;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101000;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101001;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101010;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101011;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101100;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101101;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101110;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110101111;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110000;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110001;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110010;
addr = 32'b00000000000000000101010101101110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001110110011;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110100;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110101;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110110;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110110111;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111000;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111001;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111010;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111011;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111100;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111101;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111110;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001110111111;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000000;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000001;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000010;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000011;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000100;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000101;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000110;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111000111;
addr = 32'b00000000000000000101001110110001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001111001000;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001001;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001010;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001011;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001100;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001101;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001110;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111001111;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010000;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010001;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010010;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010011;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010100;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010101;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010110;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111010111;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011000;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011001;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011010;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011011;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011100;
addr = 32'b00000000000000000101000111110100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001111011101;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011110;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111011111;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100000;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100001;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100010;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100011;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100100;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100101;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100110;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111100111;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101000;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101001;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101010;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101011;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101100;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101101;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101110;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111101111;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110000;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110001;
addr = 32'b00000000000000000101000000110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000001111110010;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110011;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110100;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110101;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110110;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111110111;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111000;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111001;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111010;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111011;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111100;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111101;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111110;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000001111111111;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000000;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000001;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000010;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000011;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000100;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000101;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000000110;
addr = 32'b00000000000000000100111001111010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010000000111;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001000;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001001;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001010;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001011;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001100;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001101;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001110;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000001111;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010000;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010001;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010010;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010011;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010100;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010101;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010110;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000010111;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011000;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011001;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011010;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011011;
addr = 32'b00000000000000000100110010111101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010000011100;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011101;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011110;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000011111;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100000;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100001;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100010;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100011;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100100;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100101;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100110;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000100111;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101000;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101001;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101010;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101011;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101100;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101101;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101110;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000101111;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110000;
addr = 32'b00000000000000000111000111011110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010000110001;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110010;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110011;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110100;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110101;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110110;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000110111;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111000;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111001;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111010;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111011;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111100;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111101;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111110;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010000111111;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000000;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000001;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000010;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000011;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000100;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000101;
addr = 32'b00000000000000000110111110111101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010001000110;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001000111;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001000;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001001;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001010;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001011;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001100;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001101;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001110;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001001111;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010000;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010001;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010010;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010011;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010100;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010101;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010110;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001010111;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011000;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011001;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011010;
addr = 32'b00000000000000000110110110011100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010001011011;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011100;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011101;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011110;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001011111;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100000;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100001;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100010;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100011;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100100;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100101;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100110;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001100111;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101000;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101001;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101010;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101011;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101100;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101101;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101110;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001101111;
addr = 32'b00000000000000000110101101111011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010001110000;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110001;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110010;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110011;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110100;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110101;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110110;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001110111;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111000;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111001;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111010;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111011;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111100;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111101;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111110;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010001111111;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000000;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000001;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000010;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000011;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000100;
addr = 32'b00000000000000000110100101011010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010010000101;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000110;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010000111;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001000;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001001;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001010;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001011;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001100;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001101;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001110;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010001111;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010000;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010001;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010010;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010011;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010100;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010101;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010110;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010010111;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011000;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011001;
addr = 32'b00000000000000000110011100111001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010010011010;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011011;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011100;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011101;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011110;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010011111;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100000;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100001;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100010;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100011;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100100;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100101;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100110;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010100111;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101000;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101001;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101010;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101011;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101100;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101101;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010101110;
addr = 32'b00000000000000000110010100011000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010010101111;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110000;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110001;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110010;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110011;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110100;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110101;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110110;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010110111;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111000;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111001;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111010;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111011;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111100;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111101;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111110;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010010111111;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000000;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000001;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000010;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000011;
addr = 32'b00000000000000000110001011110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010011000100;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000101;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000110;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011000111;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001000;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001001;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001010;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001011;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001100;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001101;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001110;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011001111;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010000;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010001;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010010;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010011;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010100;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010101;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010110;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011010111;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011000;
addr = 32'b00000000000000000110000011010110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010011011001;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011010;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011011;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011100;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011101;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011110;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011011111;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100000;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100001;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100010;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100011;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100100;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100101;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100110;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011100111;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101000;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101001;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101010;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101011;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101100;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101101;
addr = 32'b00000000000000000101111010110101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010011101110;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011101111;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110000;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110001;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110010;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110011;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110100;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110101;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110110;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011110111;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111000;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111001;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111010;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111011;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111100;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111101;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111110;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010011111111;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000000;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000001;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000010;
addr = 32'b00000000000000001000011101011010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010100000011;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000100;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000101;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000110;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100000111;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001000;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001001;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001010;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001011;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001100;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001101;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001110;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100001111;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010000;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010001;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010010;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010011;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010100;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010101;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010110;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100010111;
addr = 32'b00000000000000001000010011010101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010100011000;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011001;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011010;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011011;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011100;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011101;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011110;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100011111;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100000;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100001;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100010;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100011;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100100;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100101;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100110;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100100111;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101000;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101001;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101010;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101011;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101100;
addr = 32'b00000000000000001000001001010000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010100101101;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101110;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100101111;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110000;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110001;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110010;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110011;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110100;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110101;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110110;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100110111;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111000;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111001;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111010;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111011;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111100;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111101;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111110;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010100111111;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000000;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000001;
addr = 32'b00000000000000000111111111001011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010101000010;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000011;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000100;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000101;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000110;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101000111;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001000;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001001;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001010;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001011;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001100;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001101;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001110;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101001111;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010000;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010001;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010010;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010011;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010100;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010101;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101010110;
addr = 32'b00000000000000000111110101000110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010101010111;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011000;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011001;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011010;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011011;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011100;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011101;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011110;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101011111;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100000;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100001;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100010;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100011;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100100;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100101;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100110;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101100111;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101000;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101001;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101010;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101011;
addr = 32'b00000000000000000111101011000001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010101101100;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101101;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101110;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101101111;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110000;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110001;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110010;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110011;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110100;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110101;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110110;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101110111;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111000;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111001;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111010;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111011;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111100;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111101;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111110;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010101111111;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000000;
addr = 32'b00000000000000000111100000111100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010110000001;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000010;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000011;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000100;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000101;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000110;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110000111;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001000;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001001;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001010;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001011;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001100;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001101;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001110;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110001111;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010000;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010001;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010010;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010011;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010100;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010101;
addr = 32'b00000000000000000111010110110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010110010110;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110010111;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011000;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011001;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011010;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011011;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011100;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011101;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011110;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110011111;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100000;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100001;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100010;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100011;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100100;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100101;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100110;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110100111;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101000;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101001;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101010;
addr = 32'b00000000000000000111001100110010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010110101011;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101100;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101101;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101110;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110101111;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110000;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110001;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110010;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110011;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110100;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110101;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110110;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110110111;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111000;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111001;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111010;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111011;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111100;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111101;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111110;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010110111111;
addr = 32'b00000000000000000111000010101101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010111000000;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000001;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000010;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000011;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000100;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000101;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000110;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111000111;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001000;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001001;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001010;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001011;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001100;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001101;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001110;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111001111;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010000;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010001;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010010;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010011;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010100;
addr = 32'b00000000000000001001110011010110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010111010101;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010110;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111010111;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011000;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011001;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011010;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011011;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011100;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011101;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011110;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111011111;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100000;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100001;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100010;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100011;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100100;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100101;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100110;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111100111;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101000;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101001;
addr = 32'b00000000000000001001100111101101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010111101010;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101011;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101100;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101101;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101110;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111101111;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110000;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110001;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110010;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110011;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110100;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110101;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110110;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111110111;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111000;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111001;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111010;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111011;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111100;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111101;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000010111111110;
addr = 32'b00000000000000001001011100000100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000010111111111;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000000;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000001;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000010;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000011;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000100;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000101;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000110;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000000111;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001000;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001001;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001010;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001011;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001100;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001101;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001110;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000001111;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010000;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010001;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010010;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010011;
addr = 32'b00000000000000001001010000011011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011000010100;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010101;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010110;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000010111;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011000;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011001;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011010;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011011;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011100;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011101;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011110;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000011111;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100000;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100001;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100010;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100011;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100100;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100101;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100110;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000100111;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101000;
addr = 32'b00000000000000001001000100110010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011000101001;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101010;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101011;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101100;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101101;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101110;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000101111;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110000;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110001;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110010;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110011;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110100;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110101;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110110;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000110111;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111000;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111001;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111010;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111011;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111100;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111101;
addr = 32'b00000000000000001000111001001001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011000111110;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011000111111;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000000;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000001;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000010;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000011;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000100;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000101;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000110;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001000111;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001000;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001001;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001010;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001011;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001100;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001101;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001110;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001001111;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010000;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010001;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010010;
addr = 32'b00000000000000001000101101100000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011001010011;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010100;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010101;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010110;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001010111;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011000;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011001;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011010;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011011;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011100;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011101;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011110;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001011111;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100000;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100001;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100010;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100011;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100100;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100101;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100110;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001100111;
addr = 32'b00000000000000001000100001110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011001101000;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101001;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101010;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101011;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101100;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101101;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101110;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001101111;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110000;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110001;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110010;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110011;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110100;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110101;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110110;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001110111;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111000;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111001;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111010;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111011;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111100;
addr = 32'b00000000000000001000010110001110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011001111101;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111110;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011001111111;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000000;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000001;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000010;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000011;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000100;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000101;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000110;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010000111;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001000;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001001;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001010;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001011;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001100;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001101;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001110;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010001111;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010000;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010001;
addr = 32'b00000000000000001000001010100101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011010010010;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010011;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010100;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010101;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010110;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010010111;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011000;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011001;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011010;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011011;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011100;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011101;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011110;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010011111;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100000;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100001;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100010;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100011;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100100;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100101;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010100110;
addr = 32'b00000000000000001011001001010010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011010100111;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101000;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101001;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101010;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101011;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101100;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101101;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101110;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010101111;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110000;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110001;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110010;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110011;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110100;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110101;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110110;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010110111;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111000;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111001;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111010;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111011;
addr = 32'b00000000000000001010111100000101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011010111100;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111101;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111110;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011010111111;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000000;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000001;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000010;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000011;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000100;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000101;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000110;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011000111;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001000;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001001;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001010;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001011;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001100;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001101;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001110;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011001111;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010000;
addr = 32'b00000000000000001010101110111000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011011010001;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010010;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010011;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010100;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010101;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010110;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011010111;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011000;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011001;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011010;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011011;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011100;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011101;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011110;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011011111;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100000;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100001;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100010;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100011;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100100;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100101;
addr = 32'b00000000000000001010100001101011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011011100110;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011100111;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101000;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101001;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101010;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101011;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101100;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101101;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101110;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011101111;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110000;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110001;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110010;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110011;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110100;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110101;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110110;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011110111;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111000;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111001;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111010;
addr = 32'b00000000000000001010010100011110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011011111011;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111100;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111101;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111110;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011011111111;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000000;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000001;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000010;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000011;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000100;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000101;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000110;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100000111;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001000;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001001;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001010;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001011;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001100;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001101;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001110;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100001111;
addr = 32'b00000000000000001010000111010001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011100010000;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010001;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010010;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010011;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010100;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010101;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010110;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100010111;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011000;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011001;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011010;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011011;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011100;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011101;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011110;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100011111;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100000;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100001;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100010;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100011;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100100;
addr = 32'b00000000000000001001111010000100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011100100101;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100110;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100100111;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101000;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101001;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101010;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101011;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101100;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101101;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101110;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100101111;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110000;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110001;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110010;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110011;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110100;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110101;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110110;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100110111;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111000;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111001;
addr = 32'b00000000000000001001101100110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011100111010;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111011;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111100;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111101;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111110;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011100111111;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000000;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000001;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000010;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000011;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000100;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000101;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000110;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101000111;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001000;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001001;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001010;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001011;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001100;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001101;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101001110;
addr = 32'b00000000000000001001011111101010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011101001111;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010000;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010001;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010010;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010011;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010100;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010101;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010110;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101010111;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011000;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011001;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011010;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011011;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011100;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011101;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011110;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101011111;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100000;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100001;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100010;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100011;
addr = 32'b00000000000000001001010010011101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011101100100;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100101;
addr = 32'b00000000000000000000000001100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100110;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101100111;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101000;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101001;
addr = 32'b00000000000000000000000001010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101010;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101011;
addr = 32'b00000000000000000000000001000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101100;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101101;
addr = 32'b00000000000000000000000000111100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101110;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101101111;
addr = 32'b00000000000000000000000000110010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110000;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110001;
addr = 32'b00000000000000000000000000101000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110010;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110011;
addr = 32'b00000000000000000000000000011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110100;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110101;
addr = 32'b00000000000000000000000000010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110110;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101110111;
addr = 32'b00000000000000000000000000001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111000;
addr = 32'b00000000000000001100011111001110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011101111001;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111010;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111011;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111100;
addr = 32'b00000000000000000000000001011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111101;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111110;
addr = 32'b00000000000000000000000001001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011101111111;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000000;
addr = 32'b00000000000000000000000001000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000001;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000010;
addr = 32'b00000000000000000000000000111011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000011;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000100;
addr = 32'b00000000000000000000000000110001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000101;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000110;
addr = 32'b00000000000000000000000000100111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110000111;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001000;
addr = 32'b00000000000000000000000000011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001001;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001010;
addr = 32'b00000000000000000000000000010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001011;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001100;
addr = 32'b00000000000000000000000000001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001101;
addr = 32'b00000000000000001100010000011101;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011110001110;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110001111;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010000;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010001;
addr = 32'b00000000000000000000000001011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010010;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010011;
addr = 32'b00000000000000000000000001001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010100;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010101;
addr = 32'b00000000000000000000000001000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010110;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110010111;
addr = 32'b00000000000000000000000000111010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011000;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011001;
addr = 32'b00000000000000000000000000110000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011010;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011011;
addr = 32'b00000000000000000000000000100110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011100;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011101;
addr = 32'b00000000000000000000000000011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011110;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110011111;
addr = 32'b00000000000000000000000000010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100000;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100001;
addr = 32'b00000000000000000000000000001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100010;
addr = 32'b00000000000000001100000001101100;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011110100011;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100100;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100101;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100110;
addr = 32'b00000000000000000000000001010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110100111;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101000;
addr = 32'b00000000000000000000000001001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101001;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101010;
addr = 32'b00000000000000000000000001000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101011;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101100;
addr = 32'b00000000000000000000000000111001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101101;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101110;
addr = 32'b00000000000000000000000000101111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110101111;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110000;
addr = 32'b00000000000000000000000000100101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110001;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110010;
addr = 32'b00000000000000000000000000011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110011;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110100;
addr = 32'b00000000000000000000000000010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110101;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110110;
addr = 32'b00000000000000000000000000000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110110111;
addr = 32'b00000000000000001011110010111011;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011110111000;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111001;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111010;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111011;
addr = 32'b00000000000000000000000001010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111100;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111101;
addr = 32'b00000000000000000000000001001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111110;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011110111111;
addr = 32'b00000000000000000000000001000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000000;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000001;
addr = 32'b00000000000000000000000000111000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000010;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000011;
addr = 32'b00000000000000000000000000101110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000100;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000101;
addr = 32'b00000000000000000000000000100100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000110;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111000111;
addr = 32'b00000000000000000000000000011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001000;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001001;
addr = 32'b00000000000000000000000000010000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001010;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001011;
addr = 32'b00000000000000000000000000000110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001100;
addr = 32'b00000000000000001011100100001010;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011111001101;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001110;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111001111;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010000;
addr = 32'b00000000000000000000000001010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010001;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010010;
addr = 32'b00000000000000000000000001001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010011;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010100;
addr = 32'b00000000000000000000000001000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010101;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010110;
addr = 32'b00000000000000000000000000110111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111010111;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011000;
addr = 32'b00000000000000000000000000101101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011001;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011010;
addr = 32'b00000000000000000000000000100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011011;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011100;
addr = 32'b00000000000000000000000000011001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011101;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011110;
addr = 32'b00000000000000000000000000001111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111011111;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100000;
addr = 32'b00000000000000000000000000000101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100001;
addr = 32'b00000000000000001011010101011001;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011111100010;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100011;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100100;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100101;
addr = 32'b00000000000000000000000001010100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100110;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111100111;
addr = 32'b00000000000000000000000001001010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101000;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101001;
addr = 32'b00000000000000000000000001000000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101010;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101011;
addr = 32'b00000000000000000000000000110110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101100;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101101;
addr = 32'b00000000000000000000000000101100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101110;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111101111;
addr = 32'b00000000000000000000000000100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110000;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110001;
addr = 32'b00000000000000000000000000011000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110010;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110011;
addr = 32'b00000000000000000000000000001110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110100;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110101;
addr = 32'b00000000000000000000000000000100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111110110;
addr = 32'b00000000000000001011000110101000;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000011111110111;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111000;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111001;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111010;
addr = 32'b00000000000000000000000001010011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111011;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111100;
addr = 32'b00000000000000000000000001001001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111101;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111110;
addr = 32'b00000000000000000000000000111111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000011111111111;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000000;
addr = 32'b00000000000000000000000000110101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000001;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000010;
addr = 32'b00000000000000000000000000101011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000011;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000100;
addr = 32'b00000000000000000000000000100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000101;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000110;
addr = 32'b00000000000000000000000000010111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000000111;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001000;
addr = 32'b00000000000000000000000000001101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001001;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001010;
addr = 32'b00000000000000000000000000000011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001011;
addr = 32'b00000000000000001010110111110111;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000100000001100;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001101;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001110;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000001111;
addr = 32'b00000000000000000000000001010010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010000;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010001;
addr = 32'b00000000000000000000000001001000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010010;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010011;
addr = 32'b00000000000000000000000000111110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010100;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010101;
addr = 32'b00000000000000000000000000110100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010110;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000010111;
addr = 32'b00000000000000000000000000101010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011000;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011001;
addr = 32'b00000000000000000000000000100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011010;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011011;
addr = 32'b00000000000000000000000000010110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011100;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011101;
addr = 32'b00000000000000000000000000001100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011110;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000011111;
addr = 32'b00000000000000000000000000000010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100000;
addr = 32'b00000000000000001010101001000110;
wr = 1'b1;
#1000;

data = 32'b00000000000000000000100000100001;
addr = 32'b00000000000000000000000001011010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100010;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100011;
addr = 32'b00000000000000000000000001011011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100100;
addr = 32'b00000000000000000000000001010001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100101;
addr = 32'b00000000000000000000000001011100;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100110;
addr = 32'b00000000000000000000000001000111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000100111;
addr = 32'b00000000000000000000000001011101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101000;
addr = 32'b00000000000000000000000000111101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101001;
addr = 32'b00000000000000000000000001011110;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101010;
addr = 32'b00000000000000000000000000110011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101011;
addr = 32'b00000000000000000000000001011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101100;
addr = 32'b00000000000000000000000000101001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101101;
addr = 32'b00000000000000000000000001100000;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101110;
addr = 32'b00000000000000000000000000011111;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000101111;
addr = 32'b00000000000000000000000001100001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110000;
addr = 32'b00000000000000000000000000010101;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110001;
addr = 32'b00000000000000000000000001100010;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110010;
addr = 32'b00000000000000000000000000001011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110011;
addr = 32'b00000000000000000000000001100011;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110100;
addr = 32'b00000000000000000000000000000001;
wr = 1'b0;
#1000;

data = 32'b00000000000000000000100000110101;
addr = 32'b00000000000000001010011010010101;
wr = 1'b1;
#1000;
	$finish;	
	end
	
	always #50 clk = ~clk;			
	
	always #1000
	begin		
		if (init_state == 1)
		begin
			init_state = 0;
			#900;
		end
		if (wr == 0)
		begin
		if (is_missrate)
			missrate_counter = missrate_counter + 1;
		else
			hitrate_counter = hitrate_counter + 1;
		end
	end
	
endmodule