library verilog;
use verilog.vl_types.all;
entity cache_example is
    port(
        \out\           : out    vl_logic
    );
end cache_example;
