library verilog;
use verilog.vl_types.all;
entity rate_tb is
    port(
        a               : out    vl_logic
    );
end rate_tb;
